//START_SWREG_TABLE clint
`IOB_SWREG_W(timerInterrupt, `N_CORES-1, 0)
`IOB_SWREG_W(softwareInterrupt, `N_CORES-1, 0) 
